// Outputs all x and y values between (0,0) and (640, 480) while enable = 1
// Each value is outputted on consecutive clock cycles
// x and y begin in the top left corner and progress left to right and top to bottom
module clear_screen(clk, enable, done, x, y);
	input logic clk, enable;
	output logic done;
	output logic [10:0] x, y;
	
	always_ff @(posedge clk) begin
		if (enable) begin
			if (x == 639) begin
				x <= 0;
				if (y == 479) begin
					y <= 0;
					done <= 1'b1;
				end // if (y == 479)
				else
					y <= y + 1;
			end // if (x == 639)
			else begin
				x <= x + 1;
				if (done)
					done <= 1'b0;
			end // else
		end // if (enable)
		else begin
			x <= 0; 
			y <= 0;
			done <= 0;
		end // else
	end // always_ff
endmodule // reset_manager

module clear_screen_testbench();
	logic enable, clk, done;
	logic [10:0] x, y;
	
	// set up clock
	initial begin
		clk <= 0;
		forever #(50) clk <= ~clk;
	end // initial
	
	clear_screen dut (.*);
	
	initial begin
		enable = 0; @(posedge clk);
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		enable = 1;
		for (int i = 0; i < 307205; i++)
			@(posedge clk);
			
		$stop;
	end
endmodule // reset_manager_testbench